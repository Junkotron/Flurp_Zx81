
// Parameters used in more than one file

parameter n_periphs = 4;
parameter n_periphs_log2 = 2;
   
